module Transpose(m1, m2);
  input [0:3] m1;
  output [0:3] m2;
	
  assign m2 = m1;
endmodule
